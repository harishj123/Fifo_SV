class rst_gen;
  task rst_gen();
    #5 reset_n=1'b1;
  endtask
endclass
